// $Id: $
// File name:   test.sv
// Created:     11/8/2016
// Author:      Erin Hill
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Test for butterfly block 1
module test (
	input wire [15:0] x_0,
	input wire [15:0] x_1,
	input wire twiddle,
	output reg a_0,
	output reg a_1
);

always_comb begin
	

end



endmodule 