// $Id: $
// File name:   tb_twiddle_index3.sv
// Created:     11/24/2016
// Author:      Erin Hill
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Test bench for timer version of twiddle index
